`timescale 1ns / 1ps

module mul_LUT_20(
    input   [7:0]       in,
    output  [7:0]       out
    );
    
    reg     [7:0]       _out;
    
    assign out = _out;
    
    always @(*) begin
        casex(in)

            8'b00000000 : _out = 0;
            8'b00000001 : _out = 0;
            8'b00000010 : _out = 0;
            8'b00000011 : _out = 0;
            8'b00000100 : _out = 0;
            8'b00000101 : _out = 1;
            8'b00000110 : _out = 1;
            8'b00000111 : _out = 1;
            8'b00001000 : _out = 1;
            8'b00001001 : _out = 1;
            8'b00001010 : _out = 2;
            8'b00001011 : _out = 2;
            8'b00001100 : _out = 2;
            8'b00001101 : _out = 2;
            8'b00001110 : _out = 2;
            8'b00001111 : _out = 3;
            8'b00010000 : _out = 3;
            8'b00010001 : _out = 3;
            8'b00010010 : _out = 3;
            8'b00010011 : _out = 3;
            8'b00010100 : _out = 4;
            8'b00010101 : _out = 4;
            8'b00010110 : _out = 4;
            8'b00010111 : _out = 4;
            8'b00011000 : _out = 4;
            8'b00011001 : _out = 5;
            8'b00011010 : _out = 5;
            8'b00011011 : _out = 5;
            8'b00011100 : _out = 5;
            8'b00011101 : _out = 5;
            8'b00011110 : _out = 6;
            8'b00011111 : _out = 6;
            8'b00100000 : _out = 6;
            8'b00100001 : _out = 6;
            8'b00100010 : _out = 6;
            8'b00100011 : _out = 7;
            8'b00100100 : _out = 7;
            8'b00100101 : _out = 7;
            8'b00100110 : _out = 7;
            8'b00100111 : _out = 7;
            8'b00101000 : _out = 8;
            8'b00101001 : _out = 8;
            8'b00101010 : _out = 8;
            8'b00101011 : _out = 8;
            8'b00101100 : _out = 8;
            8'b00101101 : _out = 9;
            8'b00101110 : _out = 9;
            8'b00101111 : _out = 9;
            8'b00110000 : _out = 9;
            8'b00110001 : _out = 9;
            8'b00110010 : _out = 10;
            8'b00110011 : _out = 10;
            8'b00110100 : _out = 10;
            8'b00110101 : _out = 10;
            8'b00110110 : _out = 10;
            8'b00110111 : _out = 11;
            8'b00111000 : _out = 11;
            8'b00111001 : _out = 11;
            8'b00111010 : _out = 11;
            8'b00111011 : _out = 11;
            8'b00111100 : _out = 12;
            8'b00111101 : _out = 12;
            8'b00111110 : _out = 12;
            8'b00111111 : _out = 12;
            8'b01000000 : _out = 12;
            8'b01000001 : _out = 13;
            8'b01000010 : _out = 13;
            8'b01000011 : _out = 13;
            8'b01000100 : _out = 13;
            8'b01000101 : _out = 13;
            8'b01000110 : _out = 14;
            8'b01000111 : _out = 14;
            8'b01001000 : _out = 14;
            8'b01001001 : _out = 14;
            8'b01001010 : _out = 14;
            8'b01001011 : _out = 15;
            8'b01001100 : _out = 15;
            8'b01001101 : _out = 15;
            8'b01001110 : _out = 15;
            8'b01001111 : _out = 15;
            8'b01010000 : _out = 16;
            8'b01010001 : _out = 16;
            8'b01010010 : _out = 16;
            8'b01010011 : _out = 16;
            8'b01010100 : _out = 16;
            8'b01010101 : _out = 17;
            8'b01010110 : _out = 17;
            8'b01010111 : _out = 17;
            8'b01011000 : _out = 17;
            8'b01011001 : _out = 17;
            8'b01011010 : _out = 18;
            8'b01011011 : _out = 18;
            8'b01011100 : _out = 18;
            8'b01011101 : _out = 18;
            8'b01011110 : _out = 18;
            8'b01011111 : _out = 19;
            8'b01100000 : _out = 19;
            8'b01100001 : _out = 19;
            8'b01100010 : _out = 19;
            8'b01100011 : _out = 19;
            8'b01100100 : _out = 20;
            8'b01100101 : _out = 20;
            8'b01100110 : _out = 20;
            8'b01100111 : _out = 20;
            8'b01101000 : _out = 20;
            8'b01101001 : _out = 21;
            8'b01101010 : _out = 21;
            8'b01101011 : _out = 21;
            8'b01101100 : _out = 21;
            8'b01101101 : _out = 21;
            8'b01101110 : _out = 22;
            8'b01101111 : _out = 22;
            8'b01110000 : _out = 22;
            8'b01110001 : _out = 22;
            8'b01110010 : _out = 22;
            8'b01110011 : _out = 23;
            8'b01110100 : _out = 23;
            8'b01110101 : _out = 23;
            8'b01110110 : _out = 23;
            8'b01110111 : _out = 23;
            8'b01111000 : _out = 24;
            8'b01111001 : _out = 24;
            8'b01111010 : _out = 24;
            8'b01111011 : _out = 24;
            8'b01111100 : _out = 24;
            8'b01111101 : _out = 25;
            8'b01111110 : _out = 25;
            8'b01111111 : _out = 25;
            8'b10000000 : _out = 25;
            8'b10000001 : _out = 25;
            8'b10000010 : _out = 26;
            8'b10000011 : _out = 26;
            8'b10000100 : _out = 26;
            8'b10000101 : _out = 26;
            8'b10000110 : _out = 26;
            8'b10000111 : _out = 27;
            8'b10001000 : _out = 27;
            8'b10001001 : _out = 27;
            8'b10001010 : _out = 27;
            8'b10001011 : _out = 27;
            8'b10001100 : _out = 28;
            8'b10001101 : _out = 28;
            8'b10001110 : _out = 28;
            8'b10001111 : _out = 28;
            8'b10010000 : _out = 28;
            8'b10010001 : _out = 29;
            8'b10010010 : _out = 29;
            8'b10010011 : _out = 29;
            8'b10010100 : _out = 29;
            8'b10010101 : _out = 29;
            8'b10010110 : _out = 30;
            8'b10010111 : _out = 30;
            8'b10011000 : _out = 30;
            8'b10011001 : _out = 30;
            8'b10011010 : _out = 30;
            8'b10011011 : _out = 31;
            8'b10011100 : _out = 31;
            8'b10011101 : _out = 31;
            8'b10011110 : _out = 31;
            8'b10011111 : _out = 31;
            8'b10100000 : _out = 32;
            8'b10100001 : _out = 32;
            8'b10100010 : _out = 32;
            8'b10100011 : _out = 32;
            8'b10100100 : _out = 32;
            8'b10100101 : _out = 33;
            8'b10100110 : _out = 33;
            8'b10100111 : _out = 33;
            8'b10101000 : _out = 33;
            8'b10101001 : _out = 33;
            8'b10101010 : _out = 34;
            8'b10101011 : _out = 34;
            8'b10101100 : _out = 34;
            8'b10101101 : _out = 34;
            8'b10101110 : _out = 34;
            8'b10101111 : _out = 35;
            8'b10110000 : _out = 35;
            8'b10110001 : _out = 35;
            8'b10110010 : _out = 35;
            8'b10110011 : _out = 35;
            8'b10110100 : _out = 36;
            8'b10110101 : _out = 36;
            8'b10110110 : _out = 36;
            8'b10110111 : _out = 36;
            8'b10111000 : _out = 36;
            8'b10111001 : _out = 37;
            8'b10111010 : _out = 37;
            8'b10111011 : _out = 37;
            8'b10111100 : _out = 37;
            8'b10111101 : _out = 37;
            8'b10111110 : _out = 38;
            8'b10111111 : _out = 38;
            8'b11000000 : _out = 38;
            8'b11000001 : _out = 38;
            8'b11000010 : _out = 38;
            8'b11000011 : _out = 39;
            8'b11000100 : _out = 39;
            8'b11000101 : _out = 39;
            8'b11000110 : _out = 39;
            8'b11000111 : _out = 39;
            8'b11001000 : _out = 40;
            8'b11001001 : _out = 40;
            8'b11001010 : _out = 40;
            8'b11001011 : _out = 40;
            8'b11001100 : _out = 40;
            8'b11001101 : _out = 41;
            8'b11001110 : _out = 41;
            8'b11001111 : _out = 41;
            8'b11010000 : _out = 41;
            8'b11010001 : _out = 41;
            8'b11010010 : _out = 42;
            8'b11010011 : _out = 42;
            8'b11010100 : _out = 42;
            8'b11010101 : _out = 42;
            8'b11010110 : _out = 42;
            8'b11010111 : _out = 43;
            8'b11011000 : _out = 43;
            8'b11011001 : _out = 43;
            8'b11011010 : _out = 43;
            8'b11011011 : _out = 43;
            8'b11011100 : _out = 44;
            8'b11011101 : _out = 44;
            8'b11011110 : _out = 44;
            8'b11011111 : _out = 44;
            8'b11100000 : _out = 44;
            8'b11100001 : _out = 45;
            8'b11100010 : _out = 45;
            8'b11100011 : _out = 45;
            8'b11100100 : _out = 45;
            8'b11100101 : _out = 45;
            8'b11100110 : _out = 46;
            8'b11100111 : _out = 46;
            8'b11101000 : _out = 46;
            8'b11101001 : _out = 46;
            8'b11101010 : _out = 46;
            8'b11101011 : _out = 47;
            8'b11101100 : _out = 47;
            8'b11101101 : _out = 47;
            8'b11101110 : _out = 47;
            8'b11101111 : _out = 47;
            8'b11110000 : _out = 48;
            8'b11110001 : _out = 48;
            8'b11110010 : _out = 48;
            8'b11110011 : _out = 48;
            8'b11110100 : _out = 48;
            8'b11110101 : _out = 49;
            8'b11110110 : _out = 49;
            8'b11110111 : _out = 49;
            8'b11111000 : _out = 49;
            8'b11111001 : _out = 49;
            8'b11111010 : _out = 50;
            8'b11111011 : _out = 50;
            8'b11111100 : _out = 50;
            8'b11111101 : _out = 50;
            8'b11111110 : _out = 50;
            8'b11111111 : _out = 51;


            default: _out = 51;
        
        endcase
        
    end
endmodule