`timescale 1ns / 1ps

module mul_LUT_90(
    input   [7:0]       in,
    output  [7:0]       out
    );
    
    reg     [7:0]       _out;
    
    assign out = _out;
    
    always @(*) begin
        casex(in)

            8'b00000000 : _out = 0;
            8'b00000001 : _out = 0;
            8'b00000010 : _out = 1;
            8'b00000011 : _out = 2;
            8'b00000100 : _out = 3;
            8'b00000101 : _out = 4;
            8'b00000110 : _out = 5;
            8'b00000111 : _out = 6;
            8'b00001000 : _out = 7;
            8'b00001001 : _out = 8;
            8'b00001010 : _out = 9;
            8'b00001011 : _out = 9;
            8'b00001100 : _out = 10;
            8'b00001101 : _out = 11;
            8'b00001110 : _out = 12;
            8'b00001111 : _out = 13;
            8'b00010000 : _out = 14;
            8'b00010001 : _out = 15;
            8'b00010010 : _out = 16;
            8'b00010011 : _out = 17;
            8'b00010100 : _out = 18;
            8'b00010101 : _out = 18;
            8'b00010110 : _out = 19;
            8'b00010111 : _out = 20;
            8'b00011000 : _out = 21;
            8'b00011001 : _out = 22;
            8'b00011010 : _out = 23;
            8'b00011011 : _out = 24;
            8'b00011100 : _out = 25;
            8'b00011101 : _out = 26;
            8'b00011110 : _out = 27;
            8'b00011111 : _out = 27;
            8'b00100000 : _out = 28;
            8'b00100001 : _out = 29;
            8'b00100010 : _out = 30;
            8'b00100011 : _out = 31;
            8'b00100100 : _out = 32;
            8'b00100101 : _out = 33;
            8'b00100110 : _out = 34;
            8'b00100111 : _out = 35;
            8'b00101000 : _out = 36;
            8'b00101001 : _out = 36;
            8'b00101010 : _out = 37;
            8'b00101011 : _out = 38;
            8'b00101100 : _out = 39;
            8'b00101101 : _out = 40;
            8'b00101110 : _out = 41;
            8'b00101111 : _out = 42;
            8'b00110000 : _out = 43;
            8'b00110001 : _out = 44;
            8'b00110010 : _out = 45;
            8'b00110011 : _out = 45;
            8'b00110100 : _out = 46;
            8'b00110101 : _out = 47;
            8'b00110110 : _out = 48;
            8'b00110111 : _out = 49;
            8'b00111000 : _out = 50;
            8'b00111001 : _out = 51;
            8'b00111010 : _out = 52;
            8'b00111011 : _out = 53;
            8'b00111100 : _out = 54;
            8'b00111101 : _out = 54;
            8'b00111110 : _out = 55;
            8'b00111111 : _out = 56;
            8'b01000000 : _out = 57;
            8'b01000001 : _out = 58;
            8'b01000010 : _out = 59;
            8'b01000011 : _out = 60;
            8'b01000100 : _out = 61;
            8'b01000101 : _out = 62;
            8'b01000110 : _out = 63;
            8'b01000111 : _out = 63;
            8'b01001000 : _out = 64;
            8'b01001001 : _out = 65;
            8'b01001010 : _out = 66;
            8'b01001011 : _out = 67;
            8'b01001100 : _out = 68;
            8'b01001101 : _out = 69;
            8'b01001110 : _out = 70;
            8'b01001111 : _out = 71;
            8'b01010000 : _out = 72;
            8'b01010001 : _out = 72;
            8'b01010010 : _out = 73;
            8'b01010011 : _out = 74;
            8'b01010100 : _out = 75;
            8'b01010101 : _out = 76;
            8'b01010110 : _out = 77;
            8'b01010111 : _out = 78;
            8'b01011000 : _out = 79;
            8'b01011001 : _out = 80;
            8'b01011010 : _out = 81;
            8'b01011011 : _out = 81;
            8'b01011100 : _out = 82;
            8'b01011101 : _out = 83;
            8'b01011110 : _out = 84;
            8'b01011111 : _out = 85;
            8'b01100000 : _out = 86;
            8'b01100001 : _out = 87;
            8'b01100010 : _out = 88;
            8'b01100011 : _out = 89;
            8'b01100100 : _out = 90;
            8'b01100101 : _out = 90;
            8'b01100110 : _out = 91;
            8'b01100111 : _out = 92;
            8'b01101000 : _out = 93;
            8'b01101001 : _out = 94;
            8'b01101010 : _out = 95;
            8'b01101011 : _out = 96;
            8'b01101100 : _out = 97;
            8'b01101101 : _out = 98;
            8'b01101110 : _out = 99;
            8'b01101111 : _out = 99;
            8'b01110000 : _out = 100;
            8'b01110001 : _out = 101;
            8'b01110010 : _out = 102;
            8'b01110011 : _out = 103;
            8'b01110100 : _out = 104;
            8'b01110101 : _out = 105;
            8'b01110110 : _out = 106;
            8'b01110111 : _out = 107;
            8'b01111000 : _out = 108;
            8'b01111001 : _out = 108;
            8'b01111010 : _out = 109;
            8'b01111011 : _out = 110;
            8'b01111100 : _out = 111;
            8'b01111101 : _out = 112;
            8'b01111110 : _out = 113;
            8'b01111111 : _out = 114;
            8'b10000000 : _out = 115;
            8'b10000001 : _out = 116;
            8'b10000010 : _out = 117;
            8'b10000011 : _out = 117;
            8'b10000100 : _out = 118;
            8'b10000101 : _out = 119;
            8'b10000110 : _out = 120;
            8'b10000111 : _out = 121;
            8'b10001000 : _out = 122;
            8'b10001001 : _out = 123;
            8'b10001010 : _out = 124;
            8'b10001011 : _out = 125;
            8'b10001100 : _out = 126;
            8'b10001101 : _out = 126;
            8'b10001110 : _out = 127;
            8'b10001111 : _out = 128;
            8'b10010000 : _out = 129;
            8'b10010001 : _out = 130;
            8'b10010010 : _out = 131;
            8'b10010011 : _out = 132;
            8'b10010100 : _out = 133;
            8'b10010101 : _out = 134;
            8'b10010110 : _out = 135;
            8'b10010111 : _out = 135;
            8'b10011000 : _out = 136;
            8'b10011001 : _out = 137;
            8'b10011010 : _out = 138;
            8'b10011011 : _out = 139;
            8'b10011100 : _out = 140;
            8'b10011101 : _out = 141;
            8'b10011110 : _out = 142;
            8'b10011111 : _out = 143;
            8'b10100000 : _out = 144;
            8'b10100001 : _out = 144;
            8'b10100010 : _out = 145;
            8'b10100011 : _out = 146;
            8'b10100100 : _out = 147;
            8'b10100101 : _out = 148;
            8'b10100110 : _out = 149;
            8'b10100111 : _out = 150;
            8'b10101000 : _out = 151;
            8'b10101001 : _out = 152;
            8'b10101010 : _out = 153;
            8'b10101011 : _out = 153;
            8'b10101100 : _out = 154;
            8'b10101101 : _out = 155;
            8'b10101110 : _out = 156;
            8'b10101111 : _out = 157;
            8'b10110000 : _out = 158;
            8'b10110001 : _out = 159;
            8'b10110010 : _out = 160;
            8'b10110011 : _out = 161;
            8'b10110100 : _out = 162;
            8'b10110101 : _out = 162;
            8'b10110110 : _out = 163;
            8'b10110111 : _out = 164;
            8'b10111000 : _out = 165;
            8'b10111001 : _out = 166;
            8'b10111010 : _out = 167;
            8'b10111011 : _out = 168;
            8'b10111100 : _out = 169;
            8'b10111101 : _out = 170;
            8'b10111110 : _out = 171;
            8'b10111111 : _out = 171;
            8'b11000000 : _out = 172;
            8'b11000001 : _out = 173;
            8'b11000010 : _out = 174;
            8'b11000011 : _out = 175;
            8'b11000100 : _out = 176;
            8'b11000101 : _out = 177;
            8'b11000110 : _out = 178;
            8'b11000111 : _out = 179;
            8'b11001000 : _out = 180;
            8'b11001001 : _out = 180;
            8'b11001010 : _out = 181;
            8'b11001011 : _out = 182;
            8'b11001100 : _out = 183;
            8'b11001101 : _out = 184;
            8'b11001110 : _out = 185;
            8'b11001111 : _out = 186;
            8'b11010000 : _out = 187;
            8'b11010001 : _out = 188;
            8'b11010010 : _out = 189;
            8'b11010011 : _out = 189;
            8'b11010100 : _out = 190;
            8'b11010101 : _out = 191;
            8'b11010110 : _out = 192;
            8'b11010111 : _out = 193;
            8'b11011000 : _out = 194;
            8'b11011001 : _out = 195;
            8'b11011010 : _out = 196;
            8'b11011011 : _out = 197;
            8'b11011100 : _out = 198;
            8'b11011101 : _out = 198;
            8'b11011110 : _out = 199;
            8'b11011111 : _out = 200;
            8'b11100000 : _out = 201;
            8'b11100001 : _out = 202;
            8'b11100010 : _out = 203;
            8'b11100011 : _out = 204;
            8'b11100100 : _out = 205;
            8'b11100101 : _out = 206;
            8'b11100110 : _out = 207;
            8'b11100111 : _out = 207;
            8'b11101000 : _out = 208;
            8'b11101001 : _out = 209;
            8'b11101010 : _out = 210;
            8'b11101011 : _out = 211;
            8'b11101100 : _out = 212;
            8'b11101101 : _out = 213;
            8'b11101110 : _out = 214;
            8'b11101111 : _out = 215;
            8'b11110000 : _out = 216;
            8'b11110001 : _out = 216;
            8'b11110010 : _out = 217;
            8'b11110011 : _out = 218;
            8'b11110100 : _out = 219;
            8'b11110101 : _out = 220;
            8'b11110110 : _out = 221;
            8'b11110111 : _out = 222;
            8'b11111000 : _out = 223;
            8'b11111001 : _out = 224;
            8'b11111010 : _out = 225;
            8'b11111011 : _out = 225;
            8'b11111100 : _out = 226;
            8'b11111101 : _out = 227;
            8'b11111110 : _out = 228;
            8'b11111111 : _out = 229;


            default: _out = 229;
        
        endcase
        
    end
endmodule